// this module is an interface to use the PmodJSTK
module pmodjstk (
    // inputs / outputs
);
    // logic
endmodule