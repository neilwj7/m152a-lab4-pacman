// this module is a testbench for PmodJSTK
module pmodjstk_tb (
    // inputs + outputs
);
    // logic
endmodule