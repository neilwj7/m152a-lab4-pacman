// this module communicates with the PmodJSTK
module spi_master (
    // inputs & outputs
);
    // logic
endmodule